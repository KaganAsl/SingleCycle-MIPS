module adder(a, b, out);
input [32:0] a, b;
output [32:0] out;
assign out = a + b;
endmodule
